/u/ekke/PDIC/lab3-karthikekke/apr/work/saed32sram.lef