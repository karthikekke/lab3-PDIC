/u/ekke/PDIC/lab3-karthikekke/apr/work/saed32nm_lvt_1p9m.lef