/u/ekke/PDIC/lab3-karthikekke/cadence_cap_tech/tech.lef