/u/ekke/PDIC/lab3-karthikekke/apr/work/saed32nm_hvt_1p9m.lef